//  How to use: 
//  1. Edit the songs on the Enter Song sheet.  
//  2. Select this whole worksheet, copy it, and paste it into a new file.  
//  3. Save the file as song_rom.v. 

module song_rom (
    input clk,
    input [8:0] addr,           // The address needs to be able to access the num entries
    output reg [15:0] dout
);  

    wire [15:0] memory [383:0]; // "note memory is 16 bits wide by 512 entries long"

    always @(posedge clk)                       
        dout = memory[addr];                    

   assign memory[	  0	] =	{1'b0, 6'd21, 9'd192 };	// Note: 2F
	assign memory[	  1	] =	{1'b0, 6'd24, 9'd192 };	// Note: 2G#Ab
	assign memory[	  2	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	  3	] =	{1'b0, 6'd33, 9'd96 };	// Note: 3F
	assign memory[	  4	] =	{1'b0, 6'd36, 9'd96 };	// Note: 3G#Ab
	assign memory[	  5	] =	{1'b1, 6'd0, 9'd96 };	// Note: rest
	assign memory[	  6	] =	{1'b0, 6'd29, 9'd96 };	// Note: 3C#Db
	assign memory[	  7	] =	{1'b0, 6'd33, 9'd96 };	// Note: 3F
	assign memory[	  8	] =	{1'b1, 6'd0, 9'd72 };	// Note: rest
	assign memory[	  9	] =	{1'b0, 6'd22, 9'd216 };	// Note: 2F#Gb
	assign memory[	 10	] =	{1'b0, 6'd13, 9'd216 };	// Note: 2A
	assign memory[	 11	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 12	] =	{1'b0, 6'd28, 9'd24 };	// Note: 3C
	assign memory[	 13	] =	{1'b0, 6'd31, 9'd24 };	// Note: 3D#Eb
	assign memory[	 14	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 15	] =	{1'b0, 6'd29, 9'd24 };	// Note: 3C#Db
	assign memory[	 16	] =	{1'b0, 6'd33, 9'd24 };	// Note: 3F
	assign memory[	 17	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 18	] =	{1'b0, 6'd28, 9'd168 };	// Note: 3C
	assign memory[	 19	] =	{1'b0, 6'd31, 9'd168 };	// Note: 3D#Eb
	assign memory[	 20	] =	{1'b1, 6'd0, 9'd144 };	// Note: rest
	assign memory[	 21	] =	{1'b0, 6'd21, 9'd216 };	// Note: 2F
	assign memory[	 22	] =	{1'b0, 6'd24, 9'd216 };	// Note: 2G#Ab
	assign memory[	 23	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 24	] =	{1'b0, 6'd29, 9'd24 };	// Note: 3C#Db
	assign memory[	 25	] =	{1'b0, 6'd26, 9'd24 };	// Note: 3A#Bb
	assign memory[	 26	] =	{1'b1, 6'd0, 9'd12 };	// Note: rest
	assign memory[	 27	] =	{1'b0, 6'd28, 9'd12 };	// Note: 3C
	assign memory[	 28	] =	{1'b0, 6'd31, 9'd12 };	// Note: 3D#Eb
	assign memory[	 29	] =	{1'b1, 6'd0, 9'd12 };	// Note: rest
	assign memory[	 30	] =	{1'b0, 6'd26, 9'd120 };	// Note: 3A#Bb
	assign memory[	 31	] =	{1'b0, 6'd31, 9'd12 };	// Note: 3D#Eb
	assign memory[	 32	] =	{1'b1, 6'd0, 9'd12 };	// Note: rest
	assign memory[	 33	] =	{1'b0, 6'd33, 9'd48 };	// Note: 3F
	assign memory[	 34	] =	{1'b1, 6'd0, 9'd48 };	// Note: rest
	assign memory[	 35	] =	{1'b0, 6'd31, 9'd48 };	// Note: 3D#Eb
	assign memory[	 36	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 37	] =	{1'b0, 6'd19, 9'd216 };	// Note: 2D#Eb
	assign memory[	 38	] =	{1'b0, 6'd22, 9'd216 };	// Note: 2F#Gb
	assign memory[	 39	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 40	] =	{1'b0, 6'd24, 9'd24 };	// Note: 2G#Ab
	assign memory[	 41	] =	{1'b0, 6'd28, 9'd24 };	// Note: 3C
	assign memory[	 42	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 43	] =	{1'b0, 6'd29, 9'd24 };	// Note: 3C#Db
	assign memory[	 44	] =	{1'b0, 6'd26, 9'd24 };	// Note: 3A#Bb
	assign memory[	 45	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 46	] =	{1'b0, 6'd28, 9'd96 };	// Note: C
	assign memory[	 47	] =	{1'b0, 6'd24, 9'd72 };	// Note: 2G#Ab
	assign memory[	 48	] =	{1'b1, 6'd0, 9'd72 };	// Note: rest
	assign memory[	 49	] =	{1'b0, 6'd19, 9'd144 };	// Note: 2D#Eb
	assign memory[	 50	] =	{1'b0, 6'd17, 9'd144 };	// Note: 2C#Db
	assign memory[	 51	] =	{1'b0, 6'd22, 9'd144 };	// Note: 2F#Gb
	assign memory[	 52	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 53	] =	{1'b0, 6'd26, 9'd24 };	// Note: 3A#Bb
	assign memory[	 54	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 55	] =	{1'b0, 6'd28, 9'd24 };	// Note: 3C
	assign memory[	 56	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 57	] =	{1'b0, 6'd26, 9'd24 };	// Note: 3A#Bb
	assign memory[	 58	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 59	] =	{1'b0, 6'd31, 9'd24 };	// Note: 3D#Eb
	assign memory[	 60	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 61	] =	{1'b0, 6'd26, 9'd24 };	// Note: 3A#Bb
	assign memory[	 62	] =	{1'b0, 6'd16, 9'd72 };	// Note: 2C 
	assign memory[	 63	] =	{1'b0, 6'd19, 9'd72 };	// Note: 2D#Eb
	assign memory[	 64	] =	{1'b0, 6'd22, 9'd72 };	// Note: 2F#Gb
	assign memory[	 65	] =	{1'b0, 6'd24, 9'd24 };	// Note: 2G#Ab
	assign memory[	 66	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 67	] =	{1'b0, 6'd26, 9'd24 };	// Note: 3A#Bb
	assign memory[	 68	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 69	] =	{1'b0, 6'd24, 9'd48 };	// Note: 2G#Ab
	assign memory[	 70	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 71	] =	{1'b0, 6'd14, 9'd144 };	// Note: 2A#Bb
	assign memory[	 72	] =	{1'b0, 6'd17, 9'd144 };	// Note: 2C#Db
	assign memory[	 73	] =	{1'b0, 6'd19, 9'd144 };	// Note: 2D#Eb
	assign memory[	 74	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 75	] =	{1'b0, 6'd22, 9'd24 };	// Note: 2F#Gb
	assign memory[	 76	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 77	] =	{1'b0, 6'd24, 9'd24 };	// Note: 2G#Ab
	assign memory[	 78	] =	{1'b0, 6'd22, 9'd24 };	// Note: 2F#Gb
	assign memory[	 79	] =	{1'b0, 6'd22, 9'd72 };	
	assign memory[	 80	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 81	] =	{1'b0, 6'd16, 9'd72 };	// Note: 2C
	assign memory[	 82	] =	{1'b0, 6'd12, 9'd72 };	// Note: 1G#Ab
	assign memory[	 83	] =	{1'b0, 6'd19, 9'd72 };	// Note: 2D#Eb
	assign memory[	 84	] =	{1'b0, 6'd21, 9'd96 };	// Note: 2F
	assign memory[	 85	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 86	] =	{1'b0, 6'd17, 9'd216 };	// Note: 2C#Db
	assign memory[	 87	] =	{1'b0, 6'd14, 9'd216 };	// Note: 2A#Bb
	assign memory[	 88	] =	{1'b0, 6'd24, 9'd144 };	// Note: 2G#Ab
	assign memory[	 89	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 90	] =	{1'b0, 6'd33, 9'd24 };	// Note: 3F
	assign memory[	 91	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 92	] =	{1'b0, 6'd22, 9'd24 };	// Note: 2F#Gb
	assign memory[	 93	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 94	] =	{1'b0, 6'd21, 9'd24 };	// Note: 2F
	assign memory[	 95	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 96	] =	{1'b0, 6'd26, 9'd24 };	// Note: 3A#Bb
	assign memory[	 97	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	 98	] =	{1'b0, 6'd21, 9'd24 };	// Note: 2F
	assign memory[	 99	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	100	] =	{1'b0, 6'd10, 9'd72 };	// Note: 1F#Gb
	assign memory[	101	] =	{1'b0, 6'd19, 9'd24 };	// Note: 2D#Eb
	assign memory[	102	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	103	] =	{1'b0, 6'd21, 9'd24 };	// Note: 2F
	assign memory[	104	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	105	] =	{1'b0, 6'd19, 9'd48 };	// Note: 2D#Eb
	assign memory[	106	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	107	] =	{1'b0, 6'd9, 9'd144 };	// Note: 1F
	assign memory[	108	] =	{1'b0, 6'd24, 9'd144 };	// Note: 2G#Ab
	assign memory[	109	] =	{1'b0, 6'd14, 9'd144 };	// Note: 2A#Bb
	assign memory[	110	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	111	] =	{1'b0, 6'd17, 9'd24 };	// Note: 2C#Db
	assign memory[	112	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	113	] =	{1'b0, 6'd19, 9'd24 };	// Note: 2D#Eb
	assign memory[	114	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	115	] =	{1'b0, 6'd17, 9'd24 };	// Note: 2C#Db
	assign memory[	116	] =	{1'b1, 6'd0, 9'd42 };	// Note: rest
	assign memory[	117	] =	{1'b0, 6'd7, 9'd48 };	// Note: 1D#Eb
	assign memory[	118	] =	{1'b0, 6'd10, 9'd72 };	// Note: 1F#Gb
	assign memory[	119	] =	{1'b0, 6'd16, 9'd72 };	// Note: 2C
	assign memory[	120	] =	{1'b0, 6'd12, 9'd72 };	// Note: 1G#Ab
	assign memory[	121	] =	{1'b1, 6'd0, 9'd24 };	// Note: rest
	assign memory[	122	] =	{1'b0, 6'd1, 9'd120 };	// Note: 1A
	assign memory[	123	] =	{1'b1, 6'd0, 9'd120 };	// Note: rest
	assign memory[	124	] =	{1'b1, 6'd0, 9'd0 };	// Note: rest
	assign memory[	125	] =	{1'b1, 6'd0, 9'd0 };	// Note: rest
	assign memory[	126	] =	{1'b1, 6'd0, 9'd0 };	// Note: rest
	assign memory[	127	] =	{1'b1, 6'd0, 9'd0 };	// Note: rest
	
	// Carol of the Bells
	assign memory[	128	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	129	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	130	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	131	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	132	] =	{1'b0, 6'd25, 9'd12};	// Note: 3A
	assign memory[	133	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	134	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	135	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	136	] =	{1'b0, 6'd23, 9'd12};	// Note: 2G
	assign memory[	137	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	138	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	139	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	140	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	141	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	142	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	143	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	144	] =	{1'b0, 6'd25, 9'd12};	// Note: 3A
	assign memory[	145	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	146	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	147	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	148	] =	{1'b0, 6'd23, 9'd12};	// Note: 2G
	assign memory[	149	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	150	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	151	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	152	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	153	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	154	] =	{1'b1, 6'd30, 9'd12};	// Note: 3D
	assign memory[	155	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	156	] =	{1'b0, 6'd25, 9'd12};	// Note: 3A
	assign memory[	157	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	158	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	159	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	160	] =	{1'b0, 6'd23, 9'd12};	// Note: 2G
	assign memory[	161	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	162	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	163	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	164	] =	{1'b0, 6'd50, 9'd72};	// Note: 5A#Bb
	assign memory[	165	] =	{1'b0, 6'd54, 9'd72};	// Note: 5D
	assign memory[	166	] =	{1'b0, 6'd59, 9'd72};	// Note: 5G
	assign memory[	167	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	168	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	169	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	170	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	171	] =	{1'b0, 6'd25, 9'd12};	// Note: 3A
	assign memory[	172	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	173	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	174	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	175	] =	{1'b0, 6'd23, 9'd12};	// Note: 2G
	assign memory[	176	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	177	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	178	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	179	] =	{1'b0, 6'd49, 9'd72};	// Note: 5A 
	assign memory[	180	] =	{1'b0, 6'd52, 9'd72};	// Note: 5C
	assign memory[	181	] =	{1'b0, 6'd57, 9'd72};	// Note: 5F
	assign memory[	182	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	183	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	184	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	185	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	186	] =	{1'b0, 6'd25, 9'd12};	// Note: 3A
	assign memory[	187	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	188	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	189	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	190	] =	{1'b0, 6'd23, 9'd12};	// Note: 2G
	assign memory[	191	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	192	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	193	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	194	] =	{1'b0, 6'd47, 9'd72};	// Note: 4G
	assign memory[	195	] =	{1'b0, 6'd50, 9'd72};	// Note: 5A#Bb
	assign memory[	196	] =	{1'b0, 6'd55, 9'd72};	// Note: 5D#Eb
	assign memory[	197	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	198	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	199	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	200	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	201	] =	{1'b0, 6'd25, 9'd12};	// Note: 3A
	assign memory[	202	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	203	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	204	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	205	] =	{1'b0, 6'd23, 9'd12};	// Note: 2G
	assign memory[	206	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	207	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	208	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	209	] =	{1'b0, 6'd54, 9'd72};	// Note: 5D
	assign memory[	210	] =	{1'b0, 6'd50, 9'd72};	// Note: 5A#Bb
	assign memory[	211	] =	{1'b0, 6'd47, 9'd72};	// Note: 4G 
	assign memory[	212	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	213	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	214	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	215	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	216	] =	{1'b0, 6'd25, 9'd12};	// Note: 3A
	assign memory[	217	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	218	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	219	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	220	] =	{1'b0, 6'd23, 9'd12};	// Note: 2G
	assign memory[	221	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	222	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	223	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	224	] =	{1'b0, 6'd47, 9'd72};	// Note: 4G
	assign memory[	225	] =	{1'b0, 6'd50, 9'd72};	// Note: 5A#Bb
	assign memory[	226	] =	{1'b0, 6'd55, 9'd72};	// Note: 5D#Eb
	assign memory[	227	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	228	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	229	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	230	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	231	] =	{1'b0, 6'd25, 9'd12};	// Note: 3A
	assign memory[	232	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	233	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	234	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	235	] =	{1'b0, 6'd23, 9'd12};	// Note: 2G
	assign memory[	236	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	237	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	238	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	239	] =	{1'b0, 6'd45, 9'd72};	// Note: 4F
	assign memory[	240	] =	{1'b0, 6'd50, 9'd72};	// Note: 5A#Bb
	assign memory[	241	] =	{1'b0, 6'd54, 9'd72};	// Note: 5D
	assign memory[	242	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	243	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	244	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	245	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	246	] =	{1'b0, 6'd25, 9'd12};	// Note: 3A
	assign memory[	247	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	248	] =	{1'b0, 6'd26, 9'd12};	// Note: 3A#Bb
	assign memory[	249	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	250	] =	{1'b0, 6'd23, 9'd12};	// Note: 2G
	assign memory[	251	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	252	] =	{1'b0, 6'd30, 9'd12};	// Note: 3D
	assign memory[	253	] =	{1'b1, 6'd0, 9'd12};	// Note: rest
	assign memory[	254	] =	{1'b0, 6'd42, 9'd12};	// Note: 4D
	assign memory[	255	] =	{1'b0, 6'd42, 9'd12};	// Note: 4D
		
	// POLONAISE
	assign memory[	256	] =	{1'b0, 6'd41, 9'd120};	// Note: 4C#Db
	assign memory[	257	] =	{1'b0, 6'd45, 9'd120};	// Note: 4F
	assign memory[	258	] =	{1'b0, 6'd12, 9'd20};	// Note: 1G#Ab
	assign memory[	259	] =	{1'b1, 6'd0, 9'd20};	// Note: rest
	assign memory[	260	] =	{1'b0, 6'd19, 9'd20};	// Note: 2D#E
	assign memory[	261	] =	{1'b0, 6'd31, 9'd20};	// Note: 3D#Eb
	assign memory[	262	] =	{1'b0, 6'd16, 9'd20};	// Note: 2C
	assign memory[	263	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	264	] =	{1'b0, 6'd40, 9'd5};	// Note: 4C
	assign memory[	265	] =	{1'b0, 6'd43, 9'd5};	// Note: 4D#Eb
	assign memory[	266	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	267	] =	{1'b0, 6'd40, 9'd40};	// Note: 4C
	assign memory[	268	] =	{1'b0, 6'd43, 9'd40};	// Note: 4D#Eb
	assign memory[	269	] =	{1'b0, 6'd24, 9'd20};	// Note: 2G#Ab
	assign memory[	270	] =	{1'b0, 6'd28, 9'd20};	// Note: 3C
	assign memory[	271	] =	{1'b0, 6'd36, 9'd20};	// Note: 3G#Ab
	assign memory[	272	] =	{1'b1, 6'd0, 9'd20};	// Note: rest
	assign memory[	273	] =	{1'b0, 6'd7, 9'd20};	// Note: 1D#Eb
	assign memory[	274	] =	{1'b0, 6'd19, 9'd20};	// Note: 2D#Eb
	assign memory[	275	] =	{1'b1, 6'd0, 9'd20};	// Note: rest
	assign memory[	276	] =	{1'b0, 6'd12, 9'd20};	// Note: 1G#Ab
	assign memory[	277	] =	{1'b0, 6'd24, 9'd20};	// Note: 2G#Ab
	assign memory[	278	] =	{1'b1, 6'd0, 9'd20};	// Note: rest
	assign memory[	279	] =	{1'b0, 6'd7, 9'd20};	// Note: 1D#Eb
	assign memory[	280	] =	{1'b0, 6'd36, 9'd5};	// Note: 3G#Ab
	assign memory[	281	] =	{1'b0, 6'd40, 9'd5};	// Note: 4C
	assign memory[	282	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	283	] =	{1'b0, 6'd38, 9'd5};	// Note: 4A#Bb
	assign memory[	284	] =	{1'b0, 6'd41, 9'd5};	// Note: 4C#Db
	assign memory[	285	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	286	] =	{1'b0, 6'd24, 9'd20};	// Note: 2G#Ab
	assign memory[	287	] =	{1'b0, 6'd41, 9'd5};	// Note: 4C#Db
	assign memory[	288	] =	{1'b0, 6'd45, 9'd5};	// Note: 4F
	assign memory[	289	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	290	] =	{1'b0, 6'd38, 9'd5};	// Note: 4A#Bb
	assign memory[	291	] =	{1'b0, 6'd40, 9'd5};	// Note: 4C
	assign memory[	292	] =	{1'b0, 6'd43, 9'd5};	// Note: 4D#Eb
	assign memory[	293	] =	{1'b1, 6'd0, 9'd6};	// Note: rest
	assign memory[	294	] =	{1'b0, 6'd45, 9'd2};	// Note: 4F
	assign memory[	295	] =	{1'b1, 6'd0, 9'd4};	// Note: rest
	assign memory[	296	] =	{1'b0, 6'd40, 9'd10};	// Note: 4C
	assign memory[	297	] =	{1'b0, 6'd43, 9'd10};	// Note: 4D#Eb
	assign memory[	298	] =	{1'b0, 6'd31, 9'd20};	// Note: 3D#Eb
	assign memory[	299	] =	{1'b0, 6'd19, 9'd20};	// Note: 2D#Eb
	assign memory[	300	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	301	] =	{1'b0, 6'd39, 9'd10};	// Note: 4B
	assign memory[	302	] =	{1'b0, 6'd42, 9'd10};	// Note: 4D
	assign memory[	303	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	304	] =	{1'b0, 6'd40, 9'd80};	// Note: 4C
	assign memory[	305	] =	{1'b0, 6'd43, 9'd80};	// Note: 4D#Eb
	assign memory[	306	] =	{1'b0, 6'd24, 9'd20};	// Note: 2G#Ab
	assign memory[	307	] =	{1'b0, 6'd28, 9'd20};	// Note: 3C
	assign memory[	308	] =	{1'b0, 6'd36, 9'd20};	// Note: 3G#Ab
	assign memory[	309	] =	{1'b1, 6'd0, 9'd20};	// Note: rest
	assign memory[	310	] =	{1'b0, 6'd7, 9'd20};	// Note: 1D#Eb
	assign memory[	311	] =	{1'b0, 6'd19, 9'd20};	// Note: 2D#Eb
	assign memory[	312	] =	{1'b1, 6'd0, 9'd20};	// Note: rest
	assign memory[	313	] =	{1'b0, 6'd12, 9'd20};	// Note: 1G#Ab
	assign memory[	314	] =	{1'b0, 6'd24, 9'd20};	// Note: 2G#Ab
	assign memory[	315	] =	{1'b0, 6'd0, 9'd20};	// Note: rest
	assign memory[	316	] =	{1'b1, 6'd7, 9'd20};	// Note: 1D#Eb
	assign memory[	317	] =	{1'b0, 6'd36, 9'd10};	// Note: 3G#Ab
	assign memory[	318	] =	{1'b0, 6'd40, 9'd10};	// Note: 4C
	assign memory[	319	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	320	] =	{1'b0, 6'd38, 9'd10};	// Note: 4A#Bb
	assign memory[	321	] =	{1'b0, 6'd41, 9'd10};	// Note: 4C#Db
	assign memory[	322	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	323	] =	{1'b0, 6'd41, 9'd10};	// Note: 4C#Db
	assign memory[	324	] =	{1'b0, 6'd45, 9'd10};	// Note: 4F
	assign memory[	325	] =	{1'b0, 6'd12, 9'd20};	// Note: 1G#Ab
	assign memory[	326	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	327	] =	{1'b0, 6'd40, 9'd10};	// Note: 4C
	assign memory[	328	] =	{1'b0, 6'd43, 9'd10};	// Note: 4D#Eb
	assign memory[	329	] =	{1'b1, 6'd0, 9'd6};	// Note: rest
	assign memory[	330	] =	{1'b0, 6'd45, 9'd2};	// Note: 4F
	assign memory[	331	] =	{1'b1, 6'd0, 9'd4};	// Note: rest
	assign memory[	332	] =	{1'b0, 6'd40, 9'd10};	// Note: 4C
	assign memory[	333	] =	{1'b0, 6'd43, 9'd10};	// Note: 4D#Eb
	assign memory[	334	] =	{1'b0, 6'd19, 9'd20};	// Note: 2D#Eb
	assign memory[	335	] =	{1'b0, 6'd31, 9'd20};	// Note: 3D#Eb
	assign memory[	336	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	337	] =	{1'b0, 6'd39, 9'd10};	// Note: 4B
	assign memory[	338	] =	{1'b0, 6'd42, 9'd10};	// Note: 4D
	assign memory[	339	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	340	] =	{1'b0, 6'd43, 9'd10};	// Note: 4D#Eb
	assign memory[	341	] =	{1'b0, 6'd45, 9'd10};	// Note: 4F
	assign memory[	342	] =	{1'b0, 6'd24, 9'd20};	// Note: 2G#Ab
	assign memory[	343	] =	{1'b0, 6'd28, 9'd20};	// Note: 3C
	assign memory[	344	] =	{1'b0, 6'd36, 9'd20};	// Note: 3G#Ab
	assign memory[	345	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	346	] =	{1'b0, 6'd40, 9'd10};	// Note: 4C
	assign memory[	347	] =	{1'b0, 6'd43, 9'd10};	// Note: 4D#Eb
	assign memory[	348	] =	{1'b1, 6'd0, 9'd6};	// Note: rest
	assign memory[	349	] =	{1'b0, 6'd45, 9'd2};	// Note: 4F
	assign memory[	350	] =	{1'b1, 6'd0, 9'd4};	// Note: rest
	assign memory[	351	] =	{1'b0, 6'd40, 9'd10};	// Note: 4C
	assign memory[	352	] =	{1'b0, 6'd43, 9'd10};	// Note: 4D#Eb
	assign memory[	353	] =	{1'b0, 6'd7, 9'd20};	// Note: 1D#Eb
	assign memory[	354	] =	{1'b0, 6'd19, 9'd20};	// Note: 2D#Eb
	assign memory[	355	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	356	] =	{1'b0, 6'd38, 9'd10};	// Note: 4A#Bb
	assign memory[	357	] =	{1'b0, 6'd42, 9'd10};	// Note: 4D
	assign memory[	358	] =	{1'b1, 6'd0, 9'd10};	// Note: rest
	assign memory[	359	] =	{1'b0, 6'd40, 9'd20};	// Note: 4C
	assign memory[	360	] =	{1'b0, 6'd43, 9'd20};	// Note: 4D#Eb
	assign memory[	361	] =	{1'b0, 6'd12, 9'd20};	// Note: 1G#Ab
	assign memory[	362	] =	{1'b0, 6'd24, 9'd20};	// Note: 2G#Ab
	assign memory[	363	] =	{1'b1, 6'd0, 9'd20};	// Note: rest
	assign memory[	364	] =	{1'b0, 6'd19, 9'd20};	// Note: 2D#Eb
	assign memory[	365	] =	{1'b0, 6'd14, 9'd20};	// Note: 2A#Bb
	assign memory[	366	] =	{1'b0, 6'd22, 9'd20};	// Note: 2F#Gb
	assign memory[	367	] =	{1'b0, 6'd43, 9'd20};	// Note: 4D#Eb
	assign memory[	368	] =	{1'b0, 6'd37, 9'd20};	// Note: 4A
	assign memory[	369	] =	{1'b0, 6'd46, 9'd20};	// Note: 4F#Gb
	assign memory[	370	] =	{1'b1, 6'd0, 9'd20};	// Note: rest
	assign memory[	371	] =	{1'b0, 6'd19, 9'd20};	// Note: 2D#Eb
	assign memory[	372	] =	{1'b0, 6'd37, 9'd20};	// Note: 4A
	assign memory[	373	] =	{1'b0, 6'd45, 9'd20};	// Note: 4F
	assign memory[	374	] =	{1'b0, 6'd16, 9'd20};	// Note: 2C
	assign memory[	375	] =	{1'b0, 6'd19, 9'd20};	// Note: 2D#Eb
	assign memory[	376	] =	{1'b0, 6'd25, 9'd20};	// Note: 3A
	assign memory[	377	] =	{1'b1, 6'd0, 9'd20};	// Note: rest
	assign memory[	378	] =	{1'b0, 6'd33, 9'd20};	// Note: 3F
	assign memory[	379	] =	{1'b0, 6'd36, 9'd480};	// Note: 3G#Ab
	assign memory[	380	] =	{1'b0, 6'd40, 9'd480};	// Note: 4C
	assign memory[	381	] =	{1'b0, 6'd31, 9'd480};	// Note: 3D#Eb
	assign memory[	382	] =	{1'b0, 6'd21, 9'd480};	// Note: 2F
	assign memory[	383	] =	{1'b0, 6'd24, 9'd480};	// Note: 2G#Ab
endmodule                           
